----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:20:07 06/07/2023 
-- Design Name: 
-- Module Name:    divider - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
-- Divider
entity divider is
    Port ( A : in  signed(7 downto 0);
           B : in  signed(7 downto 0);
           quotient : out  signed(7 downto 0));
end entity divider;

-- Divider
architecture behavioral of divider is
begin
    process (A, B)
    begin
        if B /= 0 then
            quotient <= A / B;
        else
            quotient <= (others => '0');
        end if;
    end process;
end architecture behavioral;